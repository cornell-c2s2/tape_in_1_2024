VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tapeins_sp24_tapein1_Interconnect
  CLASS BLOCK ;
  FOREIGN tapeins_sp24_tapein1_Interconnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END VPWR
  PIN adapter_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 2099.530 0.000 2099.810 4.000 ;
    END
  END adapter_parity
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 699.750 1756.000 700.030 1760.000 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END cs
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 34.040 2800.000 34.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 659.640 2800.000 660.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 722.200 2800.000 722.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 784.760 2800.000 785.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 847.320 2800.000 847.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 909.880 2800.000 910.480 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 972.440 2800.000 973.040 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1035.000 2800.000 1035.600 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1097.560 2800.000 1098.160 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1160.120 2800.000 1160.720 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1222.680 2800.000 1223.280 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 96.600 2800.000 97.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1285.240 2800.000 1285.840 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1347.800 2800.000 1348.400 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1410.360 2800.000 1410.960 ;
    END
  END io_oeb[22]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 159.160 2800.000 159.760 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 221.720 2800.000 222.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 284.280 2800.000 284.880 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 346.840 2800.000 347.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 409.400 2800.000 410.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 471.960 2800.000 472.560 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 534.520 2800.000 535.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 597.080 2800.000 597.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1472.920 2800.000 1473.520 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1535.480 2800.000 1536.080 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1598.040 2800.000 1598.640 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1660.600 2800.000 1661.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1723.160 2800.000 1723.760 ;
    END
  END io_out[4]
  PIN minion_parity
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END minion_parity
  PIN miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END miso
  PIN mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END mosi
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2099.530 1756.000 2099.810 1760.000 ;
    END
  END reset
  PIN sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1538.200 4.000 1538.800 ;
    END
  END sclk
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 10.640 2795.350 1749.200 ;
      LAYER met2 ;
        RECT 4.690 1755.720 699.470 1756.000 ;
        RECT 700.310 1755.720 2099.250 1756.000 ;
        RECT 2100.090 1755.720 2795.330 1756.000 ;
        RECT 4.690 4.280 2795.330 1755.720 ;
        RECT 4.690 4.000 699.470 4.280 ;
        RECT 700.310 4.000 2099.250 4.280 ;
        RECT 2100.090 4.000 2795.330 4.280 ;
      LAYER met3 ;
        RECT 4.000 1724.160 2796.000 1749.125 ;
        RECT 4.000 1722.760 2795.600 1724.160 ;
        RECT 4.000 1661.600 2796.000 1722.760 ;
        RECT 4.000 1660.200 2795.600 1661.600 ;
        RECT 4.000 1599.040 2796.000 1660.200 ;
        RECT 4.000 1597.640 2795.600 1599.040 ;
        RECT 4.000 1539.200 2796.000 1597.640 ;
        RECT 4.400 1537.800 2796.000 1539.200 ;
        RECT 4.000 1536.480 2796.000 1537.800 ;
        RECT 4.000 1535.080 2795.600 1536.480 ;
        RECT 4.000 1473.920 2796.000 1535.080 ;
        RECT 4.000 1472.520 2795.600 1473.920 ;
        RECT 4.000 1411.360 2796.000 1472.520 ;
        RECT 4.000 1409.960 2795.600 1411.360 ;
        RECT 4.000 1348.800 2796.000 1409.960 ;
        RECT 4.000 1347.400 2795.600 1348.800 ;
        RECT 4.000 1286.240 2796.000 1347.400 ;
        RECT 4.000 1284.840 2795.600 1286.240 ;
        RECT 4.000 1223.680 2796.000 1284.840 ;
        RECT 4.000 1222.280 2795.600 1223.680 ;
        RECT 4.000 1161.120 2796.000 1222.280 ;
        RECT 4.000 1159.720 2795.600 1161.120 ;
        RECT 4.000 1099.920 2796.000 1159.720 ;
        RECT 4.400 1098.560 2796.000 1099.920 ;
        RECT 4.400 1098.520 2795.600 1098.560 ;
        RECT 4.000 1097.160 2795.600 1098.520 ;
        RECT 4.000 1036.000 2796.000 1097.160 ;
        RECT 4.000 1034.600 2795.600 1036.000 ;
        RECT 4.000 973.440 2796.000 1034.600 ;
        RECT 4.000 972.040 2795.600 973.440 ;
        RECT 4.000 910.880 2796.000 972.040 ;
        RECT 4.000 909.480 2795.600 910.880 ;
        RECT 4.000 848.320 2796.000 909.480 ;
        RECT 4.000 846.920 2795.600 848.320 ;
        RECT 4.000 785.760 2796.000 846.920 ;
        RECT 4.000 784.360 2795.600 785.760 ;
        RECT 4.000 723.200 2796.000 784.360 ;
        RECT 4.000 721.800 2795.600 723.200 ;
        RECT 4.000 660.640 2796.000 721.800 ;
        RECT 4.400 659.240 2795.600 660.640 ;
        RECT 4.000 598.080 2796.000 659.240 ;
        RECT 4.000 596.680 2795.600 598.080 ;
        RECT 4.000 535.520 2796.000 596.680 ;
        RECT 4.000 534.120 2795.600 535.520 ;
        RECT 4.000 472.960 2796.000 534.120 ;
        RECT 4.000 471.560 2795.600 472.960 ;
        RECT 4.000 410.400 2796.000 471.560 ;
        RECT 4.000 409.000 2795.600 410.400 ;
        RECT 4.000 347.840 2796.000 409.000 ;
        RECT 4.000 346.440 2795.600 347.840 ;
        RECT 4.000 285.280 2796.000 346.440 ;
        RECT 4.000 283.880 2795.600 285.280 ;
        RECT 4.000 222.720 2796.000 283.880 ;
        RECT 4.000 221.360 2795.600 222.720 ;
        RECT 4.400 221.320 2795.600 221.360 ;
        RECT 4.400 219.960 2796.000 221.320 ;
        RECT 4.000 160.160 2796.000 219.960 ;
        RECT 4.000 158.760 2795.600 160.160 ;
        RECT 4.000 97.600 2796.000 158.760 ;
        RECT 4.000 96.200 2795.600 97.600 ;
        RECT 4.000 35.040 2796.000 96.200 ;
        RECT 4.000 33.640 2795.600 35.040 ;
        RECT 4.000 10.715 2796.000 33.640 ;
      LAYER met4 ;
        RECT 310.830 518.335 327.840 1747.425 ;
        RECT 330.240 518.335 404.640 1747.425 ;
        RECT 407.040 518.335 481.440 1747.425 ;
        RECT 483.840 518.335 558.240 1747.425 ;
        RECT 560.640 518.335 635.040 1747.425 ;
        RECT 637.440 518.335 711.840 1747.425 ;
        RECT 714.240 518.335 788.640 1747.425 ;
        RECT 791.040 518.335 865.440 1747.425 ;
        RECT 867.840 518.335 942.240 1747.425 ;
        RECT 944.640 518.335 1019.040 1747.425 ;
        RECT 1021.440 518.335 1095.840 1747.425 ;
        RECT 1098.240 518.335 1172.640 1747.425 ;
        RECT 1175.040 518.335 1249.440 1747.425 ;
        RECT 1251.840 518.335 1326.240 1747.425 ;
        RECT 1328.640 518.335 1403.040 1747.425 ;
        RECT 1405.440 518.335 1479.840 1747.425 ;
        RECT 1482.240 518.335 1556.640 1747.425 ;
        RECT 1559.040 518.335 1633.440 1747.425 ;
        RECT 1635.840 518.335 1710.240 1747.425 ;
        RECT 1712.640 518.335 1787.040 1747.425 ;
        RECT 1789.440 518.335 1863.840 1747.425 ;
        RECT 1866.240 518.335 1940.640 1747.425 ;
        RECT 1943.040 518.335 2017.440 1747.425 ;
        RECT 2019.840 518.335 2094.240 1747.425 ;
        RECT 2096.640 518.335 2171.040 1747.425 ;
        RECT 2173.440 518.335 2247.840 1747.425 ;
        RECT 2250.240 518.335 2324.640 1747.425 ;
        RECT 2327.040 518.335 2394.890 1747.425 ;
      LAYER met5 ;
        RECT 310.620 541.500 2395.100 1189.100 ;
  END
END tapeins_sp24_tapein1_Interconnect
END LIBRARY

