magic
tech sky130A
magscale 1 2
timestamp 1715535929
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 2128 559070 349840
<< metal2 >>
rect 139950 351200 140006 352000
rect 419906 351200 419962 352000
rect 139950 0 140006 800
rect 419906 0 419962 800
<< obsm2 >>
rect 938 351144 139894 351200
rect 140062 351144 419850 351200
rect 420018 351144 559066 351200
rect 938 856 559066 351144
rect 938 800 139894 856
rect 140062 800 419850 856
rect 420018 800 559066 856
<< metal3 >>
rect 559200 344632 560000 344752
rect 559200 332120 560000 332240
rect 559200 319608 560000 319728
rect 0 307640 800 307760
rect 559200 307096 560000 307216
rect 559200 294584 560000 294704
rect 559200 282072 560000 282192
rect 559200 269560 560000 269680
rect 559200 257048 560000 257168
rect 559200 244536 560000 244656
rect 559200 232024 560000 232144
rect 0 219784 800 219904
rect 559200 219512 560000 219632
rect 559200 207000 560000 207120
rect 559200 194488 560000 194608
rect 559200 181976 560000 182096
rect 559200 169464 560000 169584
rect 559200 156952 560000 157072
rect 559200 144440 560000 144560
rect 0 131928 800 132048
rect 559200 131928 560000 132048
rect 559200 119416 560000 119536
rect 559200 106904 560000 107024
rect 559200 94392 560000 94512
rect 559200 81880 560000 82000
rect 559200 69368 560000 69488
rect 559200 56856 560000 56976
rect 559200 44344 560000 44464
rect 0 44072 800 44192
rect 559200 31832 560000 31952
rect 559200 19320 560000 19440
rect 559200 6808 560000 6928
<< obsm3 >>
rect 800 344832 559200 349825
rect 800 344552 559120 344832
rect 800 332320 559200 344552
rect 800 332040 559120 332320
rect 800 319808 559200 332040
rect 800 319528 559120 319808
rect 800 307840 559200 319528
rect 880 307560 559200 307840
rect 800 307296 559200 307560
rect 800 307016 559120 307296
rect 800 294784 559200 307016
rect 800 294504 559120 294784
rect 800 282272 559200 294504
rect 800 281992 559120 282272
rect 800 269760 559200 281992
rect 800 269480 559120 269760
rect 800 257248 559200 269480
rect 800 256968 559120 257248
rect 800 244736 559200 256968
rect 800 244456 559120 244736
rect 800 232224 559200 244456
rect 800 231944 559120 232224
rect 800 219984 559200 231944
rect 880 219712 559200 219984
rect 880 219704 559120 219712
rect 800 219432 559120 219704
rect 800 207200 559200 219432
rect 800 206920 559120 207200
rect 800 194688 559200 206920
rect 800 194408 559120 194688
rect 800 182176 559200 194408
rect 800 181896 559120 182176
rect 800 169664 559200 181896
rect 800 169384 559120 169664
rect 800 157152 559200 169384
rect 800 156872 559120 157152
rect 800 144640 559200 156872
rect 800 144360 559120 144640
rect 800 132128 559200 144360
rect 880 131848 559120 132128
rect 800 119616 559200 131848
rect 800 119336 559120 119616
rect 800 107104 559200 119336
rect 800 106824 559120 107104
rect 800 94592 559200 106824
rect 800 94312 559120 94592
rect 800 82080 559200 94312
rect 800 81800 559120 82080
rect 800 69568 559200 81800
rect 800 69288 559120 69568
rect 800 57056 559200 69288
rect 800 56776 559120 57056
rect 800 44544 559200 56776
rect 800 44272 559120 44544
rect 880 44264 559120 44272
rect 880 43992 559200 44264
rect 800 32032 559200 43992
rect 800 31752 559120 32032
rect 800 19520 559200 31752
rect 800 19240 559120 19520
rect 800 7008 559200 19240
rect 800 6728 559120 7008
rect 800 2143 559200 6728
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 62166 103667 65568 349485
rect 66048 103667 80928 349485
rect 81408 103667 96288 349485
rect 96768 103667 111648 349485
rect 112128 103667 127008 349485
rect 127488 103667 142368 349485
rect 142848 103667 157728 349485
rect 158208 103667 173088 349485
rect 173568 103667 188448 349485
rect 188928 103667 203808 349485
rect 204288 103667 219168 349485
rect 219648 103667 234528 349485
rect 235008 103667 249888 349485
rect 250368 103667 265248 349485
rect 265728 103667 280608 349485
rect 281088 103667 295968 349485
rect 296448 103667 311328 349485
rect 311808 103667 326688 349485
rect 327168 103667 342048 349485
rect 342528 103667 357408 349485
rect 357888 103667 372768 349485
rect 373248 103667 388128 349485
rect 388608 103667 403488 349485
rect 403968 103667 418848 349485
rect 419328 103667 434208 349485
rect 434688 103667 449568 349485
rect 450048 103667 464928 349485
rect 465408 103667 478978 349485
<< obsm5 >>
rect 62124 108300 479020 237820
<< labels >>
rlabel metal4 s 19568 2128 19888 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 419906 0 419962 800 6 adapter_parity
port 3 nsew signal output
rlabel metal2 s 139950 351200 140006 352000 6 clk
port 4 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 cs
port 5 nsew signal input
rlabel metal3 s 559200 6808 560000 6928 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 559200 131928 560000 132048 6 io_oeb[10]
port 7 nsew signal output
rlabel metal3 s 559200 144440 560000 144560 6 io_oeb[11]
port 8 nsew signal output
rlabel metal3 s 559200 156952 560000 157072 6 io_oeb[12]
port 9 nsew signal output
rlabel metal3 s 559200 169464 560000 169584 6 io_oeb[13]
port 10 nsew signal output
rlabel metal3 s 559200 181976 560000 182096 6 io_oeb[14]
port 11 nsew signal output
rlabel metal3 s 559200 194488 560000 194608 6 io_oeb[15]
port 12 nsew signal output
rlabel metal3 s 559200 207000 560000 207120 6 io_oeb[16]
port 13 nsew signal output
rlabel metal3 s 559200 219512 560000 219632 6 io_oeb[17]
port 14 nsew signal output
rlabel metal3 s 559200 232024 560000 232144 6 io_oeb[18]
port 15 nsew signal output
rlabel metal3 s 559200 244536 560000 244656 6 io_oeb[19]
port 16 nsew signal output
rlabel metal3 s 559200 19320 560000 19440 6 io_oeb[1]
port 17 nsew signal output
rlabel metal3 s 559200 257048 560000 257168 6 io_oeb[20]
port 18 nsew signal output
rlabel metal3 s 559200 269560 560000 269680 6 io_oeb[21]
port 19 nsew signal output
rlabel metal3 s 559200 282072 560000 282192 6 io_oeb[22]
port 20 nsew signal output
rlabel metal3 s 559200 31832 560000 31952 6 io_oeb[2]
port 21 nsew signal output
rlabel metal3 s 559200 44344 560000 44464 6 io_oeb[3]
port 22 nsew signal output
rlabel metal3 s 559200 56856 560000 56976 6 io_oeb[4]
port 23 nsew signal output
rlabel metal3 s 559200 69368 560000 69488 6 io_oeb[5]
port 24 nsew signal output
rlabel metal3 s 559200 81880 560000 82000 6 io_oeb[6]
port 25 nsew signal output
rlabel metal3 s 559200 94392 560000 94512 6 io_oeb[7]
port 26 nsew signal output
rlabel metal3 s 559200 106904 560000 107024 6 io_oeb[8]
port 27 nsew signal output
rlabel metal3 s 559200 119416 560000 119536 6 io_oeb[9]
port 28 nsew signal output
rlabel metal3 s 559200 294584 560000 294704 6 io_out[0]
port 29 nsew signal output
rlabel metal3 s 559200 307096 560000 307216 6 io_out[1]
port 30 nsew signal output
rlabel metal3 s 559200 319608 560000 319728 6 io_out[2]
port 31 nsew signal output
rlabel metal3 s 559200 332120 560000 332240 6 io_out[3]
port 32 nsew signal output
rlabel metal3 s 559200 344632 560000 344752 6 io_out[4]
port 33 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 minion_parity
port 34 nsew signal output
rlabel metal3 s 0 219784 800 219904 6 miso
port 35 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 mosi
port 36 nsew signal input
rlabel metal2 s 419906 351200 419962 352000 6 reset
port 37 nsew signal input
rlabel metal3 s 0 307640 800 307760 6 sclk
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 173364682
string GDS_FILE /scratch/el595/tape_in_1_2024/openlane/tapeins_sp24_tapein1_Interconnect/runs/24_05_12_11_46/results/signoff/tapeins_sp24_tapein1_Interconnect.magic.gds
string GDS_START 1859924
<< end >>

